import fidl "intf/ADAS.fidl"
/*
import fidl "../../systems/amb-ford/intf/rearviewcamclient.fidl"
import fidl "../../systems/amb-ford/intf/camerainfo.fidl"
import fidl "../../systems/amb-ford/intf/bodycontroldata.fidl"
import fidl "../../systems/amb-ford/intf/enginedata.fidl"
import fidl "../../../../contracts-orinoco2/packages/genivi/intf/fidl/org/genivi/NodeStateManager/Consumer.fidl"
import fidl "../../systems/amb-ford/intf/actvparkassist.fidl"
import fidl "../../systems/amb-ford/intf/visualparkassist.fidl"
import fidl "../../telematics/assistcall/intf/EACall.fidl"
import fidl "../../systems/illuminationctrl/intf/CIlluminationCtrl.fidl"
 */
package ADAS{

	component ADAS{
		provides interface com.harman.ADAS.AVMService as AVMInstance
		provides interface com.harman.ADAS.PASService as PASInstance
		provides interface com.harman.ADAS.ADASDiagnosis as ADASDiagInstance

		/*
		consumes interface org.harman.ford.rearviewcamclient instance dynamic as  AMB_RVCInfo
		consumes interface org.harman.ford.camerainfo instance dynamic as AMB_CameraInfo
		consumes interface org.harman.ford.bodycontroldata instance dynamic as AMB_BodyControlInfo
		consumes interface org.harman.ford.enginedata instance dynamic as AMB_EngineDataInfo
		consumes interface org.genivi.NodeStateManager.Consumer instance dynamic as NSM_ProxyInfo
		consumes interface org.harman.ford.actvparkassist instance dynamic as AMB_APAProxyInfo
		consumes interface org.harman.ford.visualparkassist instance dynamic as AMB_VPAInfo
		consumes interface com.harman.assistcall.EACall instance dynamic as assistcall_EACall
		consumes interface com.harman.voice.CIlluminationCtrl instance dynamic as Illumn_ProxyInfo
		*/
	}
}

